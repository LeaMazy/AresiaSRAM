-- Projet de stage ING4 : RISC-V
-- ECE Paris / ARESIA
-- BOOTLOADER VHDL

-- LIBRARIES
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ENTITY
entity Bootloader is
	port (
		--INPUTS
		clk 			: in std_logic;
		CS 			: in std_logic; 							--chip select
		addrInstBoot: in std_logic_vector(11 downto 0); --addr of boot instruction
		--OUTPUT
		instBoot: out std_logic_vector(31 downto 0)    --output boot instruction 
	);
end entity;

-- ARCHITECTURE
architecture archi of Bootloader is
	TYPE ROM IS ARRAY(0 TO 204) OF std_logic_vector(31 DOWNTO 0);
	SIGNAL rom_block : ROM :=(
		x"37110000",
		x"ef00c016",
		x"73001000",
		x"6f000000",
		x"130101ff",
		x"130505fe",
		x"a3070100",
		x"1375f50f",
		x"9307f003",
		x"63e2a714",
		x"93070023",
		x"13152500",
		x"3305f500",
		x"83270500",
		x"67800700",
		x"930790ff",
		x"a307f100",
		x"0345f100",
		x"13010101",
		x"67800000",
		x"930700fb",
		x"6ff0dffe",
		x"930790f9",
		x"6ff05ffe",
		x"930720f8",
		x"6ff0dffd",
		x"930780ff",
		x"6ff05ffd",
		x"930700f8",
		x"6ff0dffc",
		x"930700f9",
		x"6ff05ffc",
		x"930780f8",
		x"6ff0dffb",
		x"930730f8",
		x"6ff05ffb",
		x"930760fc",
		x"6ff0dffa",
		x"930710fa",
		x"6ff05ffa",
		x"930760f8",
		x"6ff0dff9",
		x"9307e0f8",
		x"6ff05ff9",
		x"930720fc",
		x"6ff0dff8",
		x"9307b0f8",
		x"6ff05ff8",
		x"9307b0ff",
		x"6ff0dff7",
		x"930710fe",
		x"6ff05ff7",
		x"9307a0f8",
		x"6ff0dff6",
		x"930770fc",
		x"6ff05ff6",
		x"9307a0fa",
		x"6ff0dff5",
		x"9307b0fa",
		x"6ff05ff5",
		x"930700fc",
		x"6ff0dff4",
		x"9307c0f8",
		x"6ff05ff4",
		x"930780f9",
		x"6ff0dff3",
		x"9307e0fc",
		x"6ff05ff3",
		x"930720f9",
		x"6ff0dff2",
		x"930770f8",
		x"6ff05ff2",
		x"930730fc",
		x"6ff0dff1",
		x"930750fb",
		x"6ff05ff1",
		x"930750f9",
		x"6ff0dff0",
		x"930790f8",
		x"6ff05ff0",
		x"930710f9",
		x"6ff0dfef",
		x"930740fa",
		x"6ff05fef",
		x"9307f0ff",
		x"6ff0dfee",
		x"9307f0fb",
		x"6ff05fee",
		x"930770ff",
		x"6ff0dfed",
		x"9307f007",
		x"6ff05fed",
		x"130101fe",
		x"232a9100",
		x"93074000",
		x"232c8100",
		x"232e1100",
		x"2324f100",
		x"13040000",
		x"93040033",
		x"83278100",
		x"636af406",
		x"b7070080",
		x"23a40700",
		x"23a20700",
		x"0347c100",
		x"13178700",
		x"23a4e700",
		x"0347d100",
		x"83a68700",
		x"3367d700",
		x"23a4e700",
		x"0347e100",
		x"13178701",
		x"23a2e700",
		x"0347f100",
		x"83a64700",
		x"13170701",
		x"3367d700",
		x"23a2e700",
		x"03470101",
		x"83a64700",
		x"13178700",
		x"3367d700",
		x"23a2e700",
		x"03471101",
		x"83a64700",
		x"3367d700",
		x"23a2e700",
		x"6f000000",
		x"b3079400",
		x"03c50700",
		x"eff01fe0",
		x"93070401",
		x"1375f50f",
		x"b3872700",
		x"13041400",
		x"238ea7fe",
		x"1374f40f",
		x"6ff05ff6",
		x"50010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"58010000",
		x"68010000",
		x"68010000",
		x"f0000000",
		x"3c000000",
		x"48010000",
		x"50000000",
		x"58000000",
		x"10010000",
		x"60000000",
		x"68000000",
		x"70000000",
		x"78000000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"80000000",
		x"88000000",
		x"90000000",
		x"98000000",
		x"a0000000",
		x"a8000000",
		x"b0000000",
		x"b8000000",
		x"c0000000",
		x"c8000000",
		x"d0000000",
		x"d8000000",
		x"e0000000",
		x"e8000000",
		x"f0000000",
		x"f8000000",
		x"00010000",
		x"08010000",
		x"10010000",
		x"18010000",
		x"20010000",
		x"28010000",
		x"30010000",
		x"38010000",
		x"40010000",
		x"48010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"68010000",
		x"60010000",
		x"424f4f54"
	);
	begin
	instBoot <= rom_block(to_integer(unsigned(addrInstBoot))) when (rising_edge(clk));
	
end archi;
-- END FILE