-- Projet de stage ING4 : RISC-V
-- ECE Paris / ARESIA
-- BOOTLOADER VHDL

-- LIBRARIES
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- ENTITY
entity Bootloader is
	port (
		--INPUTS
		BootClock 			: in std_logic;
		CS 					: in std_logic; 							--chip select
		BootReset			: in std_logic;
		BootStore			: in std_logic;
		BootLoad				: in std_logic;
		BootAddr				: in std_logic_vector(11 downto 0); --addr of boot instruction
		BootIn				: in std_logic_vector(31 downto 0);
		BootFunct3			: in std_logic_vector(2 downto 0);
		--OUTPUT
		BootOut				: out std_logic_vector(31 downto 0) --output boot instruction 
	);
end entity;

-- ARCHITECTURE
architecture archi of Bootloader is
	TYPE ROM IS ARRAY(0 TO 1023) OF std_logic_vector(0 to 31);
	SIGNAL rom_block : ROM :=(
		x"00001137" , x"16c000ef" , x"00100073" , x"0000006f" , x"ff010113" , x"fe050513" , x"000107a3" , x"0ff57513",
		x"03f00793" , x"14a7e263" , x"23400793" , x"00251513" , x"00f50533" , x"00052783" , x"00078067" , x"ff900793",
		x"00f107a3" , x"00f14503" , x"01010113" , x"00008067" , x"fb000793" , x"fedff06f" , x"f9900793" , x"fe5ff06f",
		x"f8200793" , x"fddff06f" , x"ff800793" , x"fd5ff06f" , x"f8000793" , x"fcdff06f" , x"f9000793" , x"fc5ff06f",
		x"f8800793" , x"fbdff06f" , x"f8300793" , x"fb5ff06f" , x"fc600793" , x"fadff06f" , x"fa100793" , x"fa5ff06f",
		x"f8600793" , x"f9dff06f" , x"f8e00793" , x"f95ff06f" , x"fc200793" , x"f8dff06f" , x"f8b00793" , x"f85ff06f",
		x"ffb00793" , x"f7dff06f" , x"fe100793" , x"f75ff06f" , x"f8a00793" , x"f6dff06f" , x"fc700793" , x"f65ff06f",
		x"faa00793" , x"f5dff06f" , x"fab00793" , x"f55ff06f" , x"fc000793" , x"f4dff06f" , x"f8c00793" , x"f45ff06f",
		x"f9800793" , x"f3dff06f" , x"fce00793" , x"f35ff06f" , x"f9200793" , x"f2dff06f" , x"f8700793" , x"f25ff06f",
		x"fc300793" , x"f1dff06f" , x"fb500793" , x"f15ff06f" , x"f9500793" , x"f0dff06f" , x"f8900793" , x"f05ff06f",
		x"f9100793" , x"efdff06f" , x"fa400793" , x"ef5ff06f" , x"fff00793" , x"eedff06f" , x"fbf00793" , x"ee5ff06f",
		x"ff700793" , x"eddff06f" , x"07f00793" , x"ed5ff06f" , x"fe010113" , x"00912a23" , x"00400793" , x"00812c23",
		x"00112e23" , x"00f12423" , x"00000413" , x"33400493" , x"00812783" , x"06f46c63" , x"00008737" , x"800007b7",
		x"3c070713" , x"00e7a423" , x"00c14703" , x"00871713" , x"00e7a423" , x"00d14703" , x"0087a683" , x"00d76733",
		x"00e7a423" , x"00e14703" , x"01871713" , x"00e7a223" , x"00f14703" , x"0047a683" , x"01071713" , x"00d76733",
		x"00e7a223" , x"01014703" , x"0047a683" , x"00871713" , x"00d76733" , x"00e7a223" , x"01114703" , x"0047a683",
		x"00d76733" , x"00e7a223" , x"0000006f" , x"009407b3" , x"0007c503" , x"dfdff0ef" , x"01040793" , x"0ff57513",
		x"002787b3" , x"00140413" , x"fea78e23" , x"0ff47413" , x"f61ff06f" , x"00000150" , x"00000168" , x"00000168",
		x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168",
		x"00000168" , x"00000168" , x"00000158" , x"00000168" , x"00000168" , x"000000f0" , x"0000003c" , x"00000148",
		x"00000050" , x"00000058" , x"00000110" , x"00000060" , x"00000068" , x"00000070" , x"00000078" , x"00000168",
		x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000080" , x"00000088",
		x"00000090" , x"00000098" , x"000000a0" , x"000000a8" , x"000000b0" , x"000000b8" , x"000000c0" , x"000000c8",
		x"000000d0" , x"000000d8" , x"000000e0" , x"000000e8" , x"000000f0" , x"000000f8" , x"00000100" , x"00000108",
		x"00000110" , x"00000118" , x"00000120" , x"00000128" , x"00000130" , x"00000138" , x"00000140" , x"00000148",
		x"00000168" , x"00000168" , x"00000168" , x"00000168" , x"00000160" , x"544f4f42" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000",
		x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" , x"00000000" 
	);
--	signal sigad : integer;
--	signal sigpc : std_logic_vector(11 downto 0);
--	begin
--		sigpc <= addrInstBoot(11 downto 0);
--		instBoot <= rom_block(sigad) when rising_edge(clk);
--		sigad <= 206 when ((unsigned(sigpc) > 1023)) else to_integer(unsigned(sigpc));
	--	instBoot <= rom_block(to_integer(unsigned(addrInstBoot))) when (rising_edge(clk));
	
	signal SigBootAddr00 : integer;
	signal SigBootAddr08 : integer;
	signal SigBootAddr16 : integer;
	signal SigBootAddr24 : integer;
	signal SigBootOut00 : std_logic_vector(31 downto 0);
	signal SigBootOut08 : std_logic_vector(31 downto 0);
	signal SigBootOut16 : std_logic_vector(31 downto 0);
	signal SigBootOut24 : std_logic_vector(31 downto 0);
	signal sigad : integer;
	signal sigpc : std_logic_vector(11 downto 0);
	
--	signal intAddr : std_logic_vector(13 downto 0);
	
	begin
	-- BEGIN
	
--	intAddr <= DMaddr(13 downto 0);
--	cs <= not DMaddr(31);
	
	-- useful adresses used to store or load
	SigBootAddr00 <= to_integer(unsigned(BootAddr)) when (CS='1' and (BootLoad = '1' OR BootStore = '1')) else
						0;
	SigBootAddr08 <= to_integer(unsigned(BootAddr)) + 1 when (CS='1' and (BootLoad = '1' OR BootStore = '1')) else
						0;
	SigBootAddr16 <= to_integer(unsigned(BootAddr)) + 2 when (CS='1' and (BootLoad = '1' OR BootStore = '1')) else
						0;
	SigBootAddr24 <= to_integer(unsigned(BootAddr)) + 3 when (CS='1' and (BootLoad = '1' OR BootStore = '1')) else
						0;
						
	-- store for synchronous data memory
	p2 : process(BootClock, BootReset)
	begin
		if(rising_edge(BootClock)) then
			if(BootStore = '1' and CS='1') then
				if(BootFunct3 = "010") then 		--SW
					rom_block(SigBootAddr00) <= BootIn(31 downto 0);
				elsif(BootFunct3 = "001") then	--SH
					rom_block(SigBootAddr00) <= "000000" & BootIn(7 downto 0);
					rom_block(SigBootAddr08) <= "000000" & BootIn(15 downto 8);
					
				elsif(BootFunct3 = "000") then	--SB
					rom_block(SigBootAddr00) <= "000000" & BootIn(7 downto 0);
					rom_block(SigBootAddr08) <= "000000" & BootIn(15 downto 8);
					rom_block(SigBootAddr16) <= "000000" & BootIn(23 downto 16);
					rom_block(SigBootAddr24) <= "000000" & BootIn(31 downto 24);
				end if;
			end if;
		end if;
	end process;
	
	-- load for asynchronous data memory
	SigBootOut00 <= (rom_block(SigBootAddr00)) when (BootLoad = '1' and SigBootAddr00<16383) else
								(others => '0');
								
	SigBootOut08 <= rom_block(SigBootAddr08) when (BootLoad = '1' AND (BootFunct3 = "001" OR BootFunct3 = "010" OR BootFunct3 = "101") and SigBootAddr00<16383) else
								(others => '1') when ( SigBootAddr00<16383 and BootLoad = '1' AND (BootFunct3 = "000" AND ((rom_block(SigBootAddr00) AND "10000000") = "10000000"))) else
								(others => '0');
	
	SigBootOut16 <=rom_block(SigBootAddr16) when (SigBootAddr00<16383 and BootLoad = '1' AND (BootFunct3 = "010")) else
								(others => '1') when (SigBootAddr00<16383 and BootLoad = '1' AND ((BootFunct3 = "000" AND ((rom_block(SigBootAddr00) AND "10000000") = "10000000")) OR (BootFunct3 = "001" AND ((rom_block(SigBootAddr08) AND "10000000") = "10000000")))) else
								(others => '0');
	
	SigBootOut24 <=rom_block(SigBootAddr24) when (SigBootAddr00<16383 and BootLoad = '1' AND (BootFunct3 = "010")) else
								(others => '1') when (SigBootAddr00<16383 and BootLoad = '1' AND ((BootFunct3 = "000" AND ((rom_block(SigBootAddr00) AND "10000000") = "10000000")) OR (BootFunct3 = "001" AND ((rom_block(SigBootAddr08) AND "10000000") = "10000000")))) else
								(others => '0');
	
	
	sigad <= 1023 when ((unsigned(BootAddr) > 1023)) else to_integer(unsigned(BootAddr));
	BootOut <= SigBootOut24(7 downto 0) & SigBootOut16(7 downto 0) & SigBootOut08(7 downto 0) & SigBootOut00(7 downto 0) when (BootLoad = '1' OR BootStore = '1') else
				  rom_block(sigad) when rising_edge(BootClock);
	-- END
	
end archi;
-- END FILE